--        ---------------------------------------
--        --     Power Smart Control | JRF | 2018

--        --            testbench
--        ---------------------------------------
     
        
--        library ieee;
--        use ieee.std_logic_1164.all;
--        use ieee.numeric_std.all;
        
--        entity tb is            
--        end tb;
        
--        architecture tb_1 of tb is
        
--            component Test_normal_mode_MUX
--                Port ( 
--                       CLK       : in   STD_LOGIC;      
--                       RST       : in   STD_LOGIC;
                       
--                       --inputs
--                       mode                        :  in   STD_LOGIC;  
                       
--                       analog_output_TEST_1        :  in   STD_LOGIC_VECTOR (11 downto 0);   
--                       analog_output_TEST_2        :  in   STD_LOGIC_VECTOR (11 downto 0); 
--                       analog_output_TEST_3        :  in   STD_LOGIC_VECTOR (11 downto 0); 
--                       analog_output_TEST_4        :  in   STD_LOGIC_VECTOR (11 downto 0); 
--                       analog_output_TEST_5        :  in   STD_LOGIC_VECTOR (11 downto 0); 
--                       analog_output_TEST_6        :  in   STD_LOGIC_VECTOR (11 downto 0); 
--                       analog_output_TEST_7        :  in   STD_LOGIC_VECTOR (11 downto 0); 
--                       analog_output_TEST_8        :  in   STD_LOGIC_VECTOR (11 downto 0); 
--                       analog_output_TEST_9        :  in   STD_LOGIC_VECTOR (11 downto 0); 
--                       analog_output_TEST_10       :  in   STD_LOGIC_VECTOR (11 downto 0); 
--                       analog_output_TEST_11       :  in   STD_LOGIC_VECTOR (11 downto 0); 
--                       analog_output_TEST_12       :  in   STD_LOGIC_VECTOR (11 downto 0); 
--                       analog_output_TEST_13       :  in   STD_LOGIC_VECTOR (11 downto 0); 
--                       analog_output_TEST_14       :  in   STD_LOGIC_VECTOR (11 downto 0); 
--                       analog_output_TEST_15       :  in   STD_LOGIC_VECTOR (11 downto 0); 
--                       analog_output_TEST_16       :  in   STD_LOGIC_VECTOR (11 downto 0); 
--                       analog_output_TEST_17       :  in   STD_LOGIC_VECTOR (11 downto 0); 
--                       analog_output_TEST_18       :  in   STD_LOGIC_VECTOR (11 downto 0); 
                                                    
--                       analog_output_NORMAL_1      :  in   STD_LOGIC_VECTOR (11 downto 0);   
--                       analog_output_NORMAL_2      :  in   STD_LOGIC_VECTOR (11 downto 0); 
--                       analog_output_NORMAL_3      :  in   STD_LOGIC_VECTOR (11 downto 0); 
--                       analog_output_NORMAL_4      :  in   STD_LOGIC_VECTOR (11 downto 0); 
--                       analog_output_NORMAL_5      :  in   STD_LOGIC_VECTOR (11 downto 0); 
--                       analog_output_NORMAL_6      :  in   STD_LOGIC_VECTOR (11 downto 0); 
--                       analog_output_NORMAL_7      :  in   STD_LOGIC_VECTOR (11 downto 0); 
--                       analog_output_NORMAL_8      :  in   STD_LOGIC_VECTOR (11 downto 0); 
--                       analog_output_NORMAL_9      :  in   STD_LOGIC_VECTOR (11 downto 0); 
--                       analog_output_NORMAL_10     :  in   STD_LOGIC_VECTOR (11 downto 0); 
--                       analog_output_NORMAL_11     :  in   STD_LOGIC_VECTOR (11 downto 0); 
--                       analog_output_NORMAL_12     :  in   STD_LOGIC_VECTOR (11 downto 0); 
--                       analog_output_NORMAL_13     :  in   STD_LOGIC_VECTOR (11 downto 0); 
--                       analog_output_NORMAL_14     :  in   STD_LOGIC_VECTOR (11 downto 0); 
--                       analog_output_NORMAL_15     :  in   STD_LOGIC_VECTOR (11 downto 0); 
--                       analog_output_NORMAL_16     :  in   STD_LOGIC_VECTOR (11 downto 0); 
--                       analog_output_NORMAL_17     :  in   STD_LOGIC_VECTOR (11 downto 0); 
--                       analog_output_NORMAL_18     :  in   STD_LOGIC_VECTOR (11 downto 0);    
                                                   
--                       DigPot_output_TEST_1        :  in   STD_LOGIC_VECTOR (9 downto 0);   
--                       DigPot_output_TEST_2        :  in   STD_LOGIC_VECTOR (9 downto 0); 
--                       DigPot_output_TEST_3        :  in   STD_LOGIC_VECTOR (9 downto 0);    
--                       DigPot_output_TEST_4        :  in   STD_LOGIC_VECTOR (9 downto 0);    
                                                    
--                       DigPot_output_NORMAL_1      :  in   STD_LOGIC_VECTOR (9 downto 0);   
--                       DigPot_output_NORMAL_2      :  in   STD_LOGIC_VECTOR (9 downto 0); 
--                       DigPot_output_NORMAL_3      :  in   STD_LOGIC_VECTOR (9 downto 0);  
--                       DigPot_output_NORMAL_4      :  in   STD_LOGIC_VECTOR (9 downto 0);  
                                                
--                       Expansor_output_TEST_1      :  in   STD_LOGIC_VECTOR (7 downto 0);  
--                       Expansor_output_TEST_2      :  in   STD_LOGIC_VECTOR (7 downto 0); 
--                       Expansor_output_TEST_3      :  in   STD_LOGIC_VECTOR (7 downto 0); 
                                                    
--                       Expansor_output_NORMAL_1    :  in   STD_LOGIC_VECTOR (7 downto 0);  
--                       Expansor_output_NORMAL_2    :  in   STD_LOGIC_VECTOR (7 downto 0); 
--                       Expansor_output_NORMAL_3    :  in   STD_LOGIC_VECTOR (7 downto 0);
                       
--                       --outputs:           
--                       analog_output_1             : out   STD_LOGIC_VECTOR (11 downto 0);   
--                       analog_output_2             : out   STD_LOGIC_VECTOR (11 downto 0); 
--                       analog_output_3             : out   STD_LOGIC_VECTOR (11 downto 0); 
--                       analog_output_4             : out   STD_LOGIC_VECTOR (11 downto 0); 
--                       analog_output_5             : out   STD_LOGIC_VECTOR (11 downto 0); 
--                       analog_output_6             : out   STD_LOGIC_VECTOR (11 downto 0); 
--                       analog_output_7             : out   STD_LOGIC_VECTOR (11 downto 0); 
--                       analog_output_8             : out   STD_LOGIC_VECTOR (11 downto 0); 
--                       analog_output_9             : out   STD_LOGIC_VECTOR (11 downto 0); 
--                       analog_output_10            : out   STD_LOGIC_VECTOR (11 downto 0); 
--                       analog_output_11            : out   STD_LOGIC_VECTOR (11 downto 0); 
--                       analog_output_12            : out   STD_LOGIC_VECTOR (11 downto 0); 
--                       analog_output_13            : out   STD_LOGIC_VECTOR (11 downto 0); 
--                       analog_output_14            : out   STD_LOGIC_VECTOR (11 downto 0); 
--                       analog_output_15            : out   STD_LOGIC_VECTOR (11 downto 0); 
--                       analog_output_16            : out   STD_LOGIC_VECTOR (11 downto 0); 
--                       analog_output_17            : out   STD_LOGIC_VECTOR (11 downto 0); 
--                       analog_output_18            : out   STD_LOGIC_VECTOR (11 downto 0); 
                       
--                       DigPot_output_1             : out   STD_LOGIC_VECTOR (9 downto 0); 
--                       DigPot_output_2             : out   STD_LOGIC_VECTOR (9 downto 0); 
--                       DigPot_output_3             : out   STD_LOGIC_VECTOR (9 downto 0); 
--                       DigPot_output_4             : out   STD_LOGIC_VECTOR (9 downto 0); 
            
--                       Expansor_output_1           : out   STD_LOGIC_VECTOR (7 downto 0);   
--                       Expansor_output_2           : out   STD_LOGIC_VECTOR (7 downto 0);   
--                       Expansor_output_3           : out   STD_LOGIC_VECTOR (7 downto 0) 
--                       ); 
--            end component;
            
--           signal CLK                         :   STD_LOGIC:='0';      
--           signal RST                         :   STD_LOGIC:='0';
--           signal mode                        :   STD_LOGIC;  
--           signal analog_output_TEST_1        :   STD_LOGIC_VECTOR (11 downto 0);   
--           signal analog_output_TEST_2        :   STD_LOGIC_VECTOR (11 downto 0); 
--           signal analog_output_TEST_3        :   STD_LOGIC_VECTOR (11 downto 0); 
--           signal analog_output_TEST_4        :   STD_LOGIC_VECTOR (11 downto 0); 
--           signal analog_output_TEST_5        :   STD_LOGIC_VECTOR (11 downto 0); 
--           signal analog_output_TEST_6        :   STD_LOGIC_VECTOR (11 downto 0); 
--           signal analog_output_TEST_7        :   STD_LOGIC_VECTOR (11 downto 0); 
--           signal analog_output_TEST_8        :   STD_LOGIC_VECTOR (11 downto 0); 
--           signal analog_output_TEST_9        :   STD_LOGIC_VECTOR (11 downto 0); 
--           signal analog_output_TEST_10       :   STD_LOGIC_VECTOR (11 downto 0); 
--           signal analog_output_TEST_11       :   STD_LOGIC_VECTOR (11 downto 0); 
--           signal analog_output_TEST_12       :   STD_LOGIC_VECTOR (11 downto 0); 
--           signal analog_output_TEST_13       :   STD_LOGIC_VECTOR (11 downto 0); 
--           signal analog_output_TEST_14       :   STD_LOGIC_VECTOR (11 downto 0); 
--           signal analog_output_TEST_15       :   STD_LOGIC_VECTOR (11 downto 0); 
--           signal analog_output_TEST_16       :   STD_LOGIC_VECTOR (11 downto 0); 
--           signal analog_output_TEST_17       :   STD_LOGIC_VECTOR (11 downto 0); 
--           signal analog_output_TEST_18       :   STD_LOGIC_VECTOR (11 downto 0);                                         
--           signal analog_output_NORMAL_1      :   STD_LOGIC_VECTOR (11 downto 0);   
--           signal analog_output_NORMAL_2      :   STD_LOGIC_VECTOR (11 downto 0); 
--           signal analog_output_NORMAL_3      :   STD_LOGIC_VECTOR (11 downto 0); 
--           signal analog_output_NORMAL_4      :   STD_LOGIC_VECTOR (11 downto 0); 
--           signal analog_output_NORMAL_5      :   STD_LOGIC_VECTOR (11 downto 0); 
--           signal analog_output_NORMAL_6      :   STD_LOGIC_VECTOR (11 downto 0); 
--           signal analog_output_NORMAL_7      :   STD_LOGIC_VECTOR (11 downto 0); 
--           signal analog_output_NORMAL_8      :   STD_LOGIC_VECTOR (11 downto 0); 
--           signal analog_output_NORMAL_9      :   STD_LOGIC_VECTOR (11 downto 0); 
--           signal analog_output_NORMAL_10     :   STD_LOGIC_VECTOR (11 downto 0); 
--           signal analog_output_NORMAL_11     :   STD_LOGIC_VECTOR (11 downto 0); 
--           signal analog_output_NORMAL_12     :   STD_LOGIC_VECTOR (11 downto 0); 
--           signal analog_output_NORMAL_13     :   STD_LOGIC_VECTOR (11 downto 0); 
--           signal analog_output_NORMAL_14     :   STD_LOGIC_VECTOR (11 downto 0); 
--           signal analog_output_NORMAL_15     :   STD_LOGIC_VECTOR (11 downto 0); 
--           signal analog_output_NORMAL_16     :   STD_LOGIC_VECTOR (11 downto 0); 
--           signal analog_output_NORMAL_17     :   STD_LOGIC_VECTOR (11 downto 0); 
--           signal analog_output_NORMAL_18     :   STD_LOGIC_VECTOR (11 downto 0); 
--           signal DigPot_output_TEST_1        :   STD_LOGIC_VECTOR (9 downto 0);   
--           signal DigPot_output_TEST_2        :   STD_LOGIC_VECTOR (9 downto 0); 
--           signal DigPot_output_TEST_3        :   STD_LOGIC_VECTOR (9 downto 0);    
--           signal DigPot_output_TEST_4        :   STD_LOGIC_VECTOR (9 downto 0);    
--           signal DigPot_output_NORMAL_1      :   STD_LOGIC_VECTOR (9 downto 0);   
--           signal DigPot_output_NORMAL_2      :   STD_LOGIC_VECTOR (9 downto 0); 
--           signal DigPot_output_NORMAL_3      :   STD_LOGIC_VECTOR (9 downto 0);  
--           signal DigPot_output_NORMAL_4      :   STD_LOGIC_VECTOR (9 downto 0);
--           signal Expansor_output_TEST_1      :   STD_LOGIC_VECTOR (7 downto 0);  
--           signal Expansor_output_TEST_2      :   STD_LOGIC_VECTOR (7 downto 0); 
--           signal Expansor_output_TEST_3      :   STD_LOGIC_VECTOR (7 downto 0); 
--           signal Expansor_output_NORMAL_1    :   STD_LOGIC_VECTOR (7 downto 0);  
--           signal Expansor_output_NORMAL_2    :   STD_LOGIC_VECTOR (7 downto 0); 
--           signal Expansor_output_NORMAL_3    :   STD_LOGIC_VECTOR (7 downto 0);
--           signal analog_output_1             :   STD_LOGIC_VECTOR (11 downto 0);   
--           signal analog_output_2             :   STD_LOGIC_VECTOR (11 downto 0); 
--           signal analog_output_3             :   STD_LOGIC_VECTOR (11 downto 0); 
--           signal analog_output_4             :   STD_LOGIC_VECTOR (11 downto 0); 
--           signal analog_output_5             :   STD_LOGIC_VECTOR (11 downto 0); 
--           signal analog_output_6             :   STD_LOGIC_VECTOR (11 downto 0); 
--           signal analog_output_7             :   STD_LOGIC_VECTOR (11 downto 0); 
--           signal analog_output_8             :   STD_LOGIC_VECTOR (11 downto 0); 
--           signal analog_output_9             :   STD_LOGIC_VECTOR (11 downto 0); 
--           signal analog_output_10            :   STD_LOGIC_VECTOR (11 downto 0); 
--           signal analog_output_11            :   STD_LOGIC_VECTOR (11 downto 0); 
--           signal analog_output_12            :   STD_LOGIC_VECTOR (11 downto 0); 
--           signal analog_output_13            :   STD_LOGIC_VECTOR (11 downto 0); 
--           signal analog_output_14            :   STD_LOGIC_VECTOR (11 downto 0); 
--           signal analog_output_15            :   STD_LOGIC_VECTOR (11 downto 0); 
--           signal analog_output_16            :   STD_LOGIC_VECTOR (11 downto 0); 
--           signal analog_output_17            :   STD_LOGIC_VECTOR (11 downto 0); 
--           signal analog_output_18            :   STD_LOGIC_VECTOR (11 downto 0); 
--           signal DigPot_output_1             :   STD_LOGIC_VECTOR (9 downto 0); 
--           signal DigPot_output_2             :   STD_LOGIC_VECTOR (9 downto 0); 
--           signal DigPot_output_3             :   STD_LOGIC_VECTOR (9 downto 0); 
--           signal DigPot_output_4             :   STD_LOGIC_VECTOR (9 downto 0);
--           signal Expansor_output_1           :   STD_LOGIC_VECTOR (7 downto 0);   
--           signal Expansor_output_2           :   STD_LOGIC_VECTOR (7 downto 0);   
--           signal Expansor_output_3           :   STD_LOGIC_VECTOR (7 downto 0);
                
--        begin
            
--            Test_normal_mode_MUX_uut: Test_normal_mode_MUX port map (
--                CLK                           => CLK                           ,
--                RST                           => RST                           ,
--                mode                          => mode                          ,
--                analog_output_TEST_1          => analog_output_TEST_1          ,
--                analog_output_TEST_2          => analog_output_TEST_2          ,
--                analog_output_TEST_3          => analog_output_TEST_3          ,
--                analog_output_TEST_4          => analog_output_TEST_4          ,
--                analog_output_TEST_5          => analog_output_TEST_5          ,
--                analog_output_TEST_6          => analog_output_TEST_6          ,
--                analog_output_TEST_7          => analog_output_TEST_7          ,
--                analog_output_TEST_8          => analog_output_TEST_8          ,
--                analog_output_TEST_9          => analog_output_TEST_9          ,
--                analog_output_TEST_10         => analog_output_TEST_10         ,
--                analog_output_TEST_11         => analog_output_TEST_11         ,
--                analog_output_TEST_12         => analog_output_TEST_12         ,
--                analog_output_TEST_13         => analog_output_TEST_13         ,
--                analog_output_TEST_14         => analog_output_TEST_14         ,
--                analog_output_TEST_15         => analog_output_TEST_15         ,
--                analog_output_TEST_16         => analog_output_TEST_16         ,
--                analog_output_TEST_17         => analog_output_TEST_17         ,
--                analog_output_TEST_18         => analog_output_TEST_18         ,
--                analog_output_NORMAL_1        => analog_output_NORMAL_1        ,
--                analog_output_NORMAL_2        => analog_output_NORMAL_2        ,
--                analog_output_NORMAL_3        => analog_output_NORMAL_3        ,
--                analog_output_NORMAL_4        => analog_output_NORMAL_4        ,
--                analog_output_NORMAL_5        => analog_output_NORMAL_5        ,
--                analog_output_NORMAL_6        => analog_output_NORMAL_6        ,
--                analog_output_NORMAL_7        => analog_output_NORMAL_7        ,
--                analog_output_NORMAL_8        => analog_output_NORMAL_8        ,
--                analog_output_NORMAL_9        => analog_output_NORMAL_9        ,
--                analog_output_NORMAL_10       => analog_output_NORMAL_10       ,
--                analog_output_NORMAL_11       => analog_output_NORMAL_11       ,
--                analog_output_NORMAL_12       => analog_output_NORMAL_12       ,
--                analog_output_NORMAL_13       => analog_output_NORMAL_13       ,
--                analog_output_NORMAL_14       => analog_output_NORMAL_14       ,
--                analog_output_NORMAL_15       => analog_output_NORMAL_15       ,
--                analog_output_NORMAL_16       => analog_output_NORMAL_16       ,
--                analog_output_NORMAL_17       => analog_output_NORMAL_17       ,
--                analog_output_NORMAL_18       => analog_output_NORMAL_18       ,
--                DigPot_output_TEST_1          => DigPot_output_TEST_1          ,
--                DigPot_output_TEST_2          => DigPot_output_TEST_2          ,
--                DigPot_output_TEST_3          => DigPot_output_TEST_3          ,
--                DigPot_output_TEST_4          => DigPot_output_TEST_4          ,
--                DigPot_output_NORMAL_1        => DigPot_output_NORMAL_1        ,
--                DigPot_output_NORMAL_2        => DigPot_output_NORMAL_2        ,
--                DigPot_output_NORMAL_3        => DigPot_output_NORMAL_3        ,
--                DigPot_output_NORMAL_4        => DigPot_output_NORMAL_4        ,
--                Expansor_output_TEST_1        => Expansor_output_TEST_1        ,
--                Expansor_output_TEST_2        => Expansor_output_TEST_2        ,
--                Expansor_output_TEST_3        => Expansor_output_TEST_3        ,
--                Expansor_output_NORMAL_1      => Expansor_output_NORMAL_1      ,
--                Expansor_output_NORMAL_2      => Expansor_output_NORMAL_2      ,
--                Expansor_output_NORMAL_3      => Expansor_output_NORMAL_3      ,
--                analog_output_1               => analog_output_1               ,
--                analog_output_2               => analog_output_2               ,
--                analog_output_3               => analog_output_3               ,
--                analog_output_4               => analog_output_4               ,
--                analog_output_5               => analog_output_5               ,
--                analog_output_6               => analog_output_6               ,
--                analog_output_7               => analog_output_7               ,
--                analog_output_8               => analog_output_8               ,
--                analog_output_9               => analog_output_9               ,
--                analog_output_10              => analog_output_10              ,
--                analog_output_11              => analog_output_11              ,
--                analog_output_12              => analog_output_12              ,
--                analog_output_13              => analog_output_13              ,
--                analog_output_14              => analog_output_14              ,
--                analog_output_15              => analog_output_15              ,
--                analog_output_16              => analog_output_16              ,
--                analog_output_17              => analog_output_17              ,
--                analog_output_18              => analog_output_18              ,
--                DigPot_output_1               => DigPot_output_1               ,
--                DigPot_output_2               => DigPot_output_2               ,
--                DigPot_output_3               => DigPot_output_3               ,
--                DigPot_output_4               => DigPot_output_4               ,
--                Expansor_output_1             => Expansor_output_1             ,
--                Expansor_output_2             => Expansor_output_2             ,
--                Expansor_output_3             => Expansor_output_3             
--            );
            
--            CLK<= not (CLK) after 5ns;
--            RST<= '0', '1' after 100 ns;
            

--            mode <='0', '1' after 1us;         
            
                         
--            analog_output_TEST_1  <= "010010111101";     
--            analog_output_TEST_2  <= "000110111101";     
--            analog_output_TEST_3  <= "011010111101";     
--            analog_output_TEST_4  <= "000000111101";     
--            analog_output_TEST_5  <= "010010111101";     
--            analog_output_TEST_6  <= "000010100001";     
--            analog_output_TEST_7  <= "000010001101";     
--            analog_output_TEST_8  <= "011110111101";     
--            analog_output_TEST_9  <= "000111111101";     
--            analog_output_TEST_10 <= "000000011101";     
--            analog_output_TEST_11 <= "000010000001";     
--            analog_output_TEST_12 <= "000110111101";     
--            analog_output_TEST_13 <= "001111111101";     
--            analog_output_TEST_14 <= "000011111101";     
--            analog_output_TEST_15 <= "000010101101";     
--            analog_output_TEST_16 <= "000010111001";     
--            analog_output_TEST_17 <= "000010011101";     
--            analog_output_TEST_18 <= "000010110001";     
--            analog_output_NORMAL_1   <= "011111000000";  
--            analog_output_NORMAL_2   <= "011111000000";  
--            analog_output_NORMAL_3   <= "011111000000";  
--            analog_output_NORMAL_4   <= "011111000000";  
--            analog_output_NORMAL_5   <= "011111000000";  
--            analog_output_NORMAL_6   <= "011111000000";  
--            analog_output_NORMAL_7   <= "011111000000";  
--            analog_output_NORMAL_8   <= "011111000000";  
--            analog_output_NORMAL_9   <= "011111000000";  
--            analog_output_NORMAL_10  <= "011111000000";  
--            analog_output_NORMAL_11  <= "011111000000";  
--            analog_output_NORMAL_12  <= "011111000000";  
--            analog_output_NORMAL_13  <= "011111000000";  
--            analog_output_NORMAL_14  <= "011111000000";  
--            analog_output_NORMAL_15  <= "011111000000";  
--            analog_output_NORMAL_16  <= "011111000000";  
--            analog_output_NORMAL_17  <= "011111000000";  
--            analog_output_NORMAL_18  <= "011111000000"; 
             
--            DigPot_output_TEST_1     <="0000111010";  
--            DigPot_output_TEST_2     <="0000111010";  
--            DigPot_output_TEST_3     <="0000111010";  
--            DigPot_output_TEST_4     <="0000111010";  
--            DigPot_output_NORMAL_1   <="0001111111";  
--            DigPot_output_NORMAL_2   <="0001111111";  
--            DigPot_output_NORMAL_3   <="0001111111";  
--            DigPot_output_NORMAL_4   <="0001111111";  
            
--            Expansor_output_TEST_1     <="10111100";
--            Expansor_output_TEST_2     <="10111100";
--            Expansor_output_TEST_3     <="10111100";
--            Expansor_output_NORMAL_1   <="10111101";
--            Expansor_output_NORMAL_2   <="10111101";
--            Expansor_output_NORMAL_3   <="10111101";
           
           
           
--        end tb_1;

